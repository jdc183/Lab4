library verilog;
use verilog.vl_types.all;
entity \_3or\ is
    port(
        \out\           : out    vl_logic;
        x               : in     vl_logic;
        y               : in     vl_logic;
        z               : in     vl_logic
    );
end \_3or\;
