library verilog;
use verilog.vl_types.all;
entity \_3and\ is
    port(
        \out\           : out    vl_logic;
        x               : in     vl_logic;
        y               : in     vl_logic;
        z               : in     vl_logic
    );
end \_3and\;
