library verilog;
use verilog.vl_types.all;
entity \_5or\ is
    port(
        \out\           : out    vl_logic;
        x               : in     vl_logic;
        y               : in     vl_logic;
        z               : in     vl_logic;
        w               : in     vl_logic;
        v               : in     vl_logic
    );
end \_5or\;
